`define SYSOPCODE 7'b1010101
`define SHAOPCODE 7'b1010100

`define systolic_addrset_FUNC 3'b000
`define systolic_calc_FUNC 3'b001

`define SHAKE_seedaddrset_FUNC 3'd0
`define SHAKE_seedset_FUNC 3'd1
`define SHAKE_squeezeonce_FUNC 3'd2
`define SHAKE_dumponce_FUNC 3'd3