`define SYSOPCODE 7'b1010101
`define systolic_addrset_FUNC 3'b000
`define systolic_calc_FUNC 3'b001